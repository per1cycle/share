// https://verilogoj.ustc.edu.cn/oj/problem/136
module top_module(
  input in, output out
);
assign out = in;
endmodule