module example1;

initial begin
    $display("hello world");
end

endmodule