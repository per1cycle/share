// https://verilogoj.ustc.edu.cn/oj/problem/30
module top_module(
  output out
);
assign out = 1;
endmodule