// https://systemverilog.dev/1.html
module example1;

initial begin
    $display("hello world");
end

endmodule