// https://verilogoj.ustc.edu.cn/oj/problem/74
module top_module( 
    input a,b,c,
    output w,x,y,z );
// 请用户在下方编辑代码
assign w = a;
assign x = b, y = b;
assign z = c;
//用户编辑到此为止
endmodule
